*CIRCUIT DE COMANDA A BECULUI
.PARAM POT1=7K
Q1 9 7 8 BC107
Q2 15 14 13 BC107
Q3 14 15 11 BC251
R4 11 10 3K
R3 10 8 1
R2 7 6 4k
R1 6 5 100
R5 12 15 {POT1}
R6 15 4 {10K-POT1}
R7 5 12 50K
R9 9 5 1
R8 3 0 4
C 11 4 0.47U
*C1 4 5 4700U
D1 4 1 D1N4007
D2 1 5 D1N4007
D3 3 5 D1N4007
D4 4 3 D1N4007
X1 5 13 4 SC10C23D
V1 1 0  SIN(0 12V 50HZ)
V2 12 4 DC 8.2V
.LIB D:\PSPICE\LIB\BC107.MOD
.LIB D:\PSPICE\LIB\BC251.MOD
.LIB D:\PSPICE\LIB\D1N4007.MOD
.LIB D:\PSPICE\LIB\SCTHYRIS.LIB
*.DC LIN V1 8 14 0.5
*.AC LIN 100 40HZ 60HZ
.TRAN 1MS 100MS
.END