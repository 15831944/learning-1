*CIRCUIT REGULATOR
.LIB
R1 1 2 100
RPOT ANOD 1 1K
C1 1 0 1U
C2 2 0 1U
X1 ANOD 2 0 2N1595
RL REDR ANOD 500
VAC 10001 10005 AC 220 SIN (0 310 50)
.model D1N4148 D Is 10E-15 Bv 1000 Rs .1
D1 10001 REDR D1N4148
D2 0 10005 D1N4148
D3 10005 REDR D1N4148
D4 0 10001 D1N4148
D5 1 ANOD D1N4148
.tran	 2.000m  .06	 0	   ; *ipsp*
.END
