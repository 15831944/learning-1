*THYRISTOR
.SUBCKT SCR 1 2 3 2 ;ANOD,CATOD,+CONTROL,-CONTROL
S1 1 5 2 6 SMOD
RG 3 4 50
VX 4 2 DC 0V
VY 5 7 DC 0V
DT 7 2 DMOD
RT 6 2 1
CT 6 2 10UF
F1 2 6 POLY(2) VX VY 0 50 11
.MODEL SMOD VSWITCH(RON=0.0125,ROFF=10E+5,VON=0.5,VOFF=0)
.MODEL DMOD D(IS=2.2E-15 BV=12V TT=0)
.ENDS SCR
